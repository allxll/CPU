`timescale 1ns/1ps

module Inst_Mem (
	input [31:0] addr,
	output [31:0] data
);

localparam ROM_SIZE = 256;
(* rom_style = "distributed" *) reg [31:0] ROMDATA[ROM_SIZE-1:0];

assign data = (addr[30:2] < ROM_SIZE)?ROMDATA[addr[30:2]]:32'b0;

integer i;
initial begin
		ROMDATA[0]  <=  32'h08000003;
		ROMDATA[1]  <=  32'h0800001f;
        ROMDATA[2]  <=  32'h08000096;
        ROMDATA[3]  <=  32'h3c084000;
        ROMDATA[4]  <=  32'h35080008;
        ROMDATA[5]  <=  32'had000000;
        ROMDATA[6]  <=  32'h3c0affff;
        ROMDATA[7]  <=  32'h354afff6;
        ROMDATA[8]  <=  32'had0afff8;
        ROMDATA[9]  <=  32'h354affff;
        ROMDATA[10] <=  32'had0afffc;
        ROMDATA[11] <=  32'h20090003;
        ROMDATA[12] <=  32'had090000;
        ROMDATA[13] <=  32'h20040003;
        ROMDATA[14] <=  32'h0c000010;
        ROMDATA[15] <=  32'h1000ffff;
        ROMDATA[16] <=  32'h23bd0008;
        ROMDATA[17] <=  32'hafbffffc;
        ROMDATA[18] <=  32'hafa40000;
        ROMDATA[19] <=  32'h28880001;
        ROMDATA[20] <=  32'h11000003;
        ROMDATA[21] <=  32'h00001026;
        ROMDATA[22] <=  32'h23bdfff8;
        ROMDATA[23] <=  32'h03e00008;
        ROMDATA[24] <=  32'h2084ffff;
        ROMDATA[25] <=  32'h0c000010;
        ROMDATA[26] <=  32'h8fa40000;
        ROMDATA[27] <=  32'h8fbffffc;
        ROMDATA[28] <=  32'h23bdfff8;
        ROMDATA[29] <=  32'h00821020;
        ROMDATA[30] <=  32'h03e00008;
        ROMDATA[31] <=  32'hafa90004;
        ROMDATA[32] <=  32'hafa80008;
        ROMDATA[33] <=  32'h00004020;
        ROMDATA[34] <=  32'h3c084000;
        ROMDATA[35] <=  32'h3129fff9;
        ROMDATA[36] <=  32'had090008;
        ROMDATA[37] <=  32'h23bd0024;
        ROMDATA[38] <=  32'hafb00000;
        ROMDATA[39] <=  32'hafa4fffc;
        ROMDATA[40] <=  32'hafa5fff8;
        ROMDATA[41] <=  32'hafaafff4;
        ROMDATA[42] <=  32'hafa2fff0;
        ROMDATA[43] <=  32'hafa3ffec;
        ROMDATA[44] <=  32'hafbfffe8;
        ROMDATA[45] <=  32'h8d100014;
        ROMDATA[46] <=  32'h00108202;
        ROMDATA[47] <=  32'h20030001;
        ROMDATA[48] <=  32'h12030006;
        ROMDATA[49] <=  32'h00031840;
        ROMDATA[50] <=  32'h12030007;
        ROMDATA[51] <=  32'h00031840;
		ROMDATA[52] <=  32'h12030008;
		ROMDATA[53] <=  32'h00031840;
		ROMDATA[54] <=  32'h12030009;
		ROMDATA[55] <=  32'h34100200;
		ROMDATA[56] <=  32'h3084000f;
		ROMDATA[57] <=  32'h08000043;
		ROMDATA[58] <=  32'h34100400;
		ROMDATA[59] <=  32'h00052102;
		ROMDATA[60] <=  32'h08000043;
		ROMDATA[61] <=  32'h34100800;
		ROMDATA[62] <=  32'h30a4000f;
		ROMDATA[63] <=  32'h08000043;
		ROMDATA[64] <=  32'h34100100;
		ROMDATA[65] <=  32'h00042102;
		ROMDATA[66] <=  32'h08000043;
		ROMDATA[67] <=  32'h0c000047;
		ROMDATA[68] <=  32'h020a8025;
		ROMDATA[69] <=  32'had100014;
		ROMDATA[70] <=  32'h08000088;
		ROMDATA[71] <=  32'h00001020;
		ROMDATA[72] <=  32'h1082001f;
		ROMDATA[73] <=  32'h20420001;
		ROMDATA[74] <=  32'h1082001f;
		ROMDATA[75] <=  32'h20420001;
		ROMDATA[76] <=  32'h1082001f;
		ROMDATA[77] <=  32'h20420001;
		ROMDATA[78] <=  32'h1082001f;
		ROMDATA[79] <=  32'h20420001;
		ROMDATA[80] <=  32'h1082001f;
        ROMDATA[81] <=  32'h20420001;
		ROMDATA[82] <=  32'h1082001f;
		ROMDATA[83] <=  32'h20420001;
		ROMDATA[84] <=  32'h1082001f;
		ROMDATA[85] <=  32'h20420001;
		ROMDATA[86] <=  32'h1082001f;
		ROMDATA[87] <=  32'h20420001;
		ROMDATA[88] <=  32'h1082001f;
		ROMDATA[89] <=  32'h20420001;
		ROMDATA[90] <=  32'h1082001f;
		ROMDATA[91] <=  32'h20420001;
		ROMDATA[92] <=  32'h1082001f;
		ROMDATA[93] <=  32'h20420001;
		ROMDATA[94] <=  32'h1082001f;
		ROMDATA[95] <=  32'h20420001;
		ROMDATA[96] <=  32'h1082001f;
		ROMDATA[97] <=  32'h20420001;
		ROMDATA[98] <=  32'h1082001f;
		ROMDATA[99] <=  32'h20420001;
		ROMDATA[100] <= 32'h1082001f;
		ROMDATA[101] <= 32'h20420001;
		ROMDATA[102] <= 32'h1082001f;
		ROMDATA[103] <= 32'h03e00008;
		ROMDATA[104] <= 32'h200a0001;
		ROMDATA[105] <= 32'h03e00008;
		ROMDATA[106] <= 32'h200a004f;
		ROMDATA[107] <= 32'h03e00008;
		ROMDATA[108] <= 32'h200a0012;
		ROMDATA[109] <= 32'h03e00008;
		ROMDATA[110] <= 32'h200a0006;
        ROMDATA[111] <= 32'h03e00008;
        ROMDATA[112] <= 32'h200a004c;
        ROMDATA[113] <= 32'h03e00008;
        ROMDATA[114] <= 32'h200a0024;
        ROMDATA[115] <= 32'h03e00008;
        ROMDATA[116] <= 32'h200a0020;
        ROMDATA[117] <= 32'h03e00008;
        ROMDATA[118] <= 32'h200a000f;
        ROMDATA[119] <= 32'h03e00008;
        ROMDATA[120] <= 32'h200a0000;
        ROMDATA[121] <= 32'h03e00008;
        ROMDATA[122] <= 32'h200a0004;
        ROMDATA[123] <= 32'h03e00008;
        ROMDATA[124] <= 32'h200a0008;
        ROMDATA[125] <= 32'h03e00008;
        ROMDATA[126] <= 32'h200a0060;
        ROMDATA[127] <= 32'h03e00008;
        ROMDATA[128] <= 32'h200a0031;
        ROMDATA[129] <= 32'h03e00008;
        ROMDATA[130] <= 32'h200a0042;
        ROMDATA[131] <= 32'h03e00008;
        ROMDATA[132] <= 32'h200a0030;
        ROMDATA[133] <= 32'h03e00008;
        ROMDATA[134] <= 32'h200a0038;
        ROMDATA[135] <= 32'h03e00008;
        ROMDATA[136] <= 32'h23bdffdc;
        ROMDATA[137] <= 32'h35290002;
        ROMDATA[138] <= 32'had090008;
        ROMDATA[139] <= 32'h8fb00000;
        ROMDATA[140] <= 32'h8fa4fffc;
        ROMDATA[141] <= 32'h8fa5fff8;
        ROMDATA[142] <= 32'h8faafff4;
        ROMDATA[143] <= 32'h8fa2fff0;
        ROMDATA[144] <= 32'h8fa3ffec;
        ROMDATA[145] <= 32'h8fbfffe8;
        ROMDATA[146] <= 32'h8fa8ffe4;
        ROMDATA[147] <= 32'h8fa9ffe0;
        ROMDATA[148] <= 32'h235afffc;
        ROMDATA[149] <= 32'h03400008;
	    for (i=150;i<ROM_SIZE;i=i+1) begin
            ROMDATA[i] <= 32'b0;
        end
end
endmodule
