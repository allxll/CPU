module testbench_ALU (
);

reg [5:0] ALUFun;
reg [31:0] A;
reg [31:0] B;
reg Sign;
wire [31:0] S;


initial begin
	$dumpfile("alu.vcd");
	$dumpvars;

	// ALUFun = 6'b000_000;   // A + B

	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 A = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 A = 2147483647;


	// ALUFun = 6'b000_001;   // A - B

	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// ALUFun = 6'b011_000;   // A & B

	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// ALUFun = 6'b011_110;    // A | B

	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;




	// ALUFun = 6'b010_110;   // A ^ B



	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;




	// ALUFun = 6'b010_001;   // ~(A|B)


	// Sign = 1;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;


	// #10 Sign = 0;
	// A = 13; B = 33;
	// #10 A = -70;
	// #10 B = 2147483647;





	// #100 ALUFun = 6'b011_010;    // A
 




	// ALUFun = 6'b100_000;    // << A[4:0]

	// Sign = 1;
	// A = 13; B = 3;
	// #10 A = -70;
	// #10 B = 27;


	// #10 Sign = 0;
	// A = 31; B = 3;
	// #10 A = -70;
	// #10 B = 27;






	// ALUFun = 6'b100_001;     // >> A[4:0] logic

	// Sign = 1;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = -70;
	// #10 B = -1;


	// #10 Sign = 1;
	// A = 31; B = 32'hf0f0_00ff;
	// #10 A = -70;
	// #10 B = -1;




	// ALUFun = 6'b100_011;    // >> A[4:0] arithmatic


	// Sign = 1;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = -70;
	// #10 B = -1;


	// #10 Sign = 1;
	// A = 31; B = 32'hf0f0_00ff;
	// #10 A = -70;
	// #10 B = -1;





	// ALUFun = 6'b110_011;    //  A == B ? 
 


	// Sign = 0;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;


	// #10 Sign = 0;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;







	// #100 ALUFun = 6'b110_001;     // A != B?



	// Sign = 0;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;


	// #10 Sign = 0;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;



	//  ALUFun = 6'b110_101;    // A < B?

	// Sign = 1;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;


	// #10 Sign = 0;
	// A = 13; B = 32'hf0f0_00ff;
	// #10 A = 32'hf0f0_00ff;
	// #10 B = 31312223;



	ALUFun = 6'b111_101;    // A <= 0?

	Sign = 1;
	A = 13; B = 32'hf0f0_00ff;
	#10 A = 32'hf0f0_00ff;
	#10 B = 31312223;


	#10 Sign = 0;
	A = 13; B = 32'hf0f0_00ff;
	#10 A = 32'hf0f0_00ff;
	#10 B = 31312223;






	#100 ALUFun = 6'b111_011;    // A < 0 ? 








	#100 ALUFun = 6'b111_111;    // A > 0 ?











	#100 $finish;
end 

ALU simple(ALUFun, A, B, Sign, S);

endmodule